// Clock gate Testbench
// ### Author : Razu Ahamed(en.razu.ahamed@gmail.com)

module tb_clk_gate;

//////////////////////////////////////////////////////////////////////////////////////////////////
//-SIGNALS
//////////////////////////////////////////////////////////////////////////////////////////////////

logic cp_i;//Clock pulse
logic e_i;//Enable
logic te_i;//Test enable
logic q_o;//Output
logic q_model;
int pass=0;
int fail=0;
//////////////////////////////////////////////////////////////////////////////////////////////////
//-RTL
//////////////////////////////////////////////////////////////////////////////////////////////////

clk_gate u_clk_gate(
  .cp_i  (cp_i),
  .e_i   (e_i ),
  .te_i  (te_i),
  .q_o   (q_o )
);

//////////////////////////////////////////////////////////////////////////////////////////////////
//-Method
//////////////////////////////////////////////////////////////////////////////////////////////////

//task start_cp_i();
//  fork
//    forever begin
//      cp_i = 1; #5;
//      cp_i = 0; #5;
//    end
//  join_none
//endtask

//////////////////////////////////////////////////////////////////////////////////////////////////
//-MODEL
//////////////////////////////////////////////////////////////////////////////////////////////////

function automatic logic q_out(logic cp_i, logic e_i, logic te_i);
logic temp;
temp = cp_i & e_i;
if(te_i==1)
  q_out =cp_i;
else
  q_out =temp;
endfunction

//////////////////////////////////////////////////////////////////////////////////////////////////
//-Procedural
//////////////////////////////////////////////////////////////////////////////////////////////////

initial
begin
  $dumpfile("dump.vcd");
  $dumpvars;
end

initial
begin
  repeat(200)
  begin
    cp_i=$urandom;
    te_i=$urandom;
    e_i =$urandom;
    q_model = q_out(cp_i,e_i,te_i);
    #2;
    if(q_o==q_model)
      pass++;
    else
      fail++;
  end
  $display("%d Time Passed",pass);
  $display("%d Time Failed",fail);
  #100 $finish;
end
endmodule
