`define DATA_IN_WIDTH 8
`define OPCODE        2
